`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:36:56 12/02/2013 
// Design Name: 
// Module Name:    get_map_address 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module get_map_address(
    input clk,
    input hcount,
    input vcount,
    input blank,
    input x,
    input y,
    output reg[11:0] addr
    );
	 
	 
	 
	 


endmodule
